library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity contador_2_bits is
   Port (clk,clr: in STD_LOGIC;
         S: out std_LOGIC_VECTOR(1 downto 0));
end contador_2_bits;

architecture ckt of contador_2_bits is

component ffjk is
   port (ck, clr, set, j, k : in  std_logic;
                          q : out std_logic);
end component;

signal FFJK1,FFJK0 :   std_logic;
signal FFJK1Q,FFJK0Q :   std_logic;
signal ENABLE , NOTCLR:   std_logic;

begin

ENABLE <= CLK;
NOTCLR <= NOT CLR;

FF0: ffJK  port map (ENABLE,NOTCLR,'1','1','1',FFJK0Q);
FF1: ffJK  port map (FFJK0,NOTCLR,'1','1','1',FFJK1Q);


FFJK1<= NOT FFJK1Q;
FFJK0<= NOT FFJK0Q;



S(1) <= FFJK1Q;
S(0) <= FFJK0Q;

end ckt;
