library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity REGISTRADOR_1_BIT is
   Port (clk,clr : in STD_LOGIC;
		E :  in STD_LOGIC;
         	S : out STD_LOGIC);
end REGISTRADOR_1_BIT;

architecture ckt of REGISTRADOR_1_BIT is

COMPONENT ffjk is
   port (ck, clr, set, j, k : in  std_logic;
                          q : out std_logic);
end COMPONENT;

signal FFJK0Q,notclr : STD_LOGIC;

begin

notclr <= not clr;
FF0: ffJK port map (clk,notclr,'1',E,'0',FFJK0Q);


S <=FFJK0Q;

end ckt;
